package wb_pkg;

  	import ncsu_pkg::*;
	`include "ncsu_macros.svh"

	`include "wb_configuration.svh"
	`include "wb_transaction.svh"
	`include "wb_transaction_random.svh"
	`include "wb_driver.svh"
	`include "wb_monitor.svh"
	`include "wb_sequence_base.svh"
	`include "wb_sequence_random.svh"
	`include "wb_agent.svh"

endpackage
