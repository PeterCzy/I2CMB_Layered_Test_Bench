package i2cmb_env_pkg;

  	import ncsu_pkg::*;
  	import i2c_pkg::*;
	import wb_pkg::*;

	`include "i2cmb_test_1.svh"

	`include "i2cmb_generator.svh"
	`include "i2cmb_predictor.svh"
	`include "i2cmb_coverage.svh"
	`include "i2cmb_env_configuration.svh"
	`include "i2cmb_scoreboard.svh"
	`include "i2cmb_environment.svh"
	`include "i2cmb_test.svh"

endpackage
