package i2c_pkg;

	import ncsu_pkg::*;
	import wb_pkg::*;

	`include "i2c_transaction.svh"
	`include "i2c_configuration.svh"
	`include "i2c_driver.svh"
	`include "i2c_monitor.svh"
	`include "i2c_agent.svh"

endpackage
